library verilog;
use verilog.vl_types.all;
entity multi_cycle_CPU_tb is
end multi_cycle_CPU_tb;
