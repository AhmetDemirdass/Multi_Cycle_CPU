library verilog;
use verilog.vl_types.all;
entity multi_cycle_CPU_vlg_vec_tst is
end multi_cycle_CPU_vlg_vec_tst;
